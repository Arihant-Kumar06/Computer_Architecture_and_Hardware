module mux8way_tb;
wire [15:0]t_out;
reg [15:0]t_a,t_b,t_c,t_d,t_e,t_f,t_g,t_h;
reg [2:0]t_sel;
mux8way my_gate(.a(t_a), .b(t_b), .c(t_c), .d(t_d), .e(t_e), .f(t_f), .g(t_g), .h(t_h), .sel(t_sel), .out(t_out));
initial begin
    $monitor("t_a=%b, t_b=%b, t_c=%b, t_d=%b, t_e=%b, t_f=%b, t_g=%b, t_h=%b, t_sel=%b, t_out=%b", t_a, t_b, t_c, t_d, t_e, t_f, t_g, t_h, t_sel, t_out);
    t_a=16'b0000000000000000;
    t_b=16'b0101010101010101;
    t_c=16'b1010101010101010;
    t_d=16'b1111111111111111;
    t_e=16'b1100110011001100;
    t_f=16'b1111000011110000;
    t_g=16'b1111111100000000;
    t_h=16'b1110001110001110;
    t_sel=000;
    #10
    t_a=16'b0000000000000000;
    t_b=16'b0101010101010101;
    t_c=16'b1010101010101010;
    t_d=16'b1111111111111111;
    t_e=16'b1100110011001100;
    t_f=16'b1111000011110000;
    t_g=16'b1111111100000000;
    t_h=16'b1110001110001110;
    t_sel=001;
    #10
    t_a=16'b0000000000000000;
    t_b=16'b0101010101010101;
    t_c=16'b1010101010101010;
    t_d=16'b1111111111111111;
    t_e=16'b1100110011001100;
    t_f=16'b1111000011110000;
    t_g=16'b1111111100000000;
    t_h=16'b1110001110001110;
    t_sel=010;
    #10
    t_a=16'b0000000000000000;
    t_b=16'b0101010101010101;
    t_c=16'b1010101010101010;
    t_d=16'b1111111111111111;
    t_e=16'b1100110011001100;
    t_f=16'b1111000011110000;
    t_g=16'b1111111100000000;
    t_h=16'b1110001110001110;
    t_sel=011;
    #10
    t_a=16'b0000000000000000;
    t_b=16'b0101010101010101;
    t_c=16'b1010101010101010;
    t_d=16'b1111111111111111;
    t_e=16'b1100110011001100;
    t_f=16'b1111000011110000;
    t_g=16'b1111111100000000;
    t_h=16'b1110001110001110;
    t_sel=100;
    #10
    t_a=16'b0000000000000000;
    t_b=16'b0101010101010101;
    t_c=16'b1010101010101010;
    t_d=16'b1111111111111111;
    t_e=16'b1100110011001100;
    t_f=16'b1111000011110000;
    t_g=16'b1111111100000000;
    t_h=16'b1110001110001110;
    t_sel=101;
    #10
    t_a=16'b0000000000000000;
    t_b=16'b0101010101010101;
    t_c=16'b1010101010101010;
    t_d=16'b1111111111111111;
    t_e=16'b1100110011001100;
    t_f=16'b1111000011110000;
    t_g=16'b1111111100000000;
    t_h=16'b1110001110001110;
    t_sel=110;
    #10
    t_a=16'b0000000000000000;
    t_b=16'b0101010101010101;
    t_c=16'b1010101010101010;
    t_d=16'b1111111111111111;
    t_e=16'b1100110011001100;
    t_f=16'b1111000011110000;
    t_g=16'b1111111100000000;
    t_h=16'b1110001110001110;
    t_sel=111;
    
end
endmodule