module notgate(x,out);
input x;
output out;
assign out=!x;
endmodule