module and16gate(
  input [15:0]x,y,
output [15:0]out
);

assign out=x&y;

endmodule